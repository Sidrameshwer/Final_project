module mul16_1(
    input [15:0] a,b,
    output [31:0] p
    );
    wire [15:0]P1;
    wire [15:0]P2;
    wire [15:0]P3;
    wire [15:0]P4;
    wire [15:1]S;
    wire [38:1]C;
    mul_8_1 m1 (a[7:0],b[7:0],P1);
    mul_8_1 m2 (a[7:0],b[15:8],P2);
    mul_8_1 m3 (a[15:8],b[7:0],P3);
    mul_8_1 m4 (a[15:8],b[15:8],P4);
    
    assign p[7:0]=P1[7:0];
    fa_df fa1 (P1[8],P2[0],P3[0],p[8],C[1]);
    fa_df fa2 (P1[9],P2[1],P3[1],S[1],C[2]);
    fa_df fa3 (P1[10],P2[2],P3[2],S[2],C[3]);
    fa_df fa4 (P1[11],P2[3],P3[3],S[3],C[4]);
    fa_df fa5 (P1[12],P2[4],P3[4],S[4],C[5]);
    fa_df fa6 (P1[13],P2[5],P3[5],S[5],C[6]);
    fa_df fa7 (P1[14],P2[6],P3[6],S[6],C[7]);
    fa_df fa8 (P1[15],P2[7],P3[7],S[7],C[8]);
    
    fa_df fa9 (P2[8],P3[8],P4[0],S[8],C[9]);
    fa_df fa10 (P2[9],P3[9],P4[1],S[9],C[10]);
    fa_df fa11 (P2[10],P3[10],P4[2],S[10],C[11]);
    fa_df fa12 (P2[11],P3[11],P4[3],S[11],C[12]);
    fa_df fa13 (P2[12],P3[12],P4[4],S[12],C[13]);
    fa_df fa14 (P2[13],P3[13],P4[5],S[13],C[14]);
    fa_df fa15 (P2[14],P3[14],P4[6],S[14],C[15]);
    fa_df fa16 (P2[15],P3[15],P4[7],S[15],C[16]);
    
    ha_df ha1(S[1],C[1],p[9],C[17]);
    fa_df fa17(S[2],C[2],C[17],p[10],C[18]);
    fa_df fa18(S[3],C[3],C[18],p[11],C[19]);
    fa_df fa19(S[4],C[4],C[19],p[12],C[20]);
    fa_df fa20(S[5],C[5],C[20],p[13],C[21]);
    fa_df fa21(S[6],C[6],C[21],p[14],C[22]);
    fa_df fa22(S[7],C[7],C[22],p[15],C[23]);
    fa_df fa23(S[8],C[8],C[23],p[16],C[24]);
    fa_df fa24(S[9],C[9],C[24],p[17],C[25]);
    fa_df fa25(S[10],C[10],C[25],p[18],C[26]);
    fa_df fa26(S[11],C[11],C[26],p[19],C[27]);
    fa_df fa27(S[12],C[12],C[27],p[20],C[28]);
    fa_df fa28(S[13],C[13],C[28],p[21],C[29]);
    fa_df fa29(S[14],C[14],C[29],p[22],C[30]);
    fa_df fa30(S[15],C[15],C[30],p[23],C[31]);
    
    fa_df fa31(P4[8],C[16],C[31],p[24],C[32]);
    ha_df ha2(P4[9],C[32],p[25],C[33]);
    ha_df ha3(P4[10],C[33],p[26],C[34]);
    ha_df ha4(P4[11],C[34],p[27],C[35]);
    ha_df ha5(P4[12],C[35],p[28],C[36]);
    ha_df ha6(P4[13],C[36],p[29],C[37]);
    ha_df ha7(P4[14],C[37],p[30],C[38]);
    xor x1(p[31],P4[15],C[38]);
endmodule
